// helper param list for interface

parameter ENV_CMD_SIZE = 4;
typedef bit [ENV_CMD_SIZE-1:0] reg_cmd_t;

parameter ENV_DATA_SIZE = 32;
typedef bit [ENV_DATA_SIZE-1:0] req_data_t;
